module suma_logica(
    input A,
    input B,
    output S

);
    assign S = A + B;
endmodule