module complemento(
    input A,
    input B,
    output S
);
    assign S = ~A; // Se niega solo A
endmodule

